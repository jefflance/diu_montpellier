<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>31.1277,-26.4051,99.9115,-70.8303</PageViewport>
<gate>
<ID>2</ID>
<type>AE_DFF_LOW</type>
<position>48,-46</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>5 </output>
<input>
<ID>clock</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4</ID>
<type>AE_DFF_LOW</type>
<position>60,-46</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>6 </output>
<input>
<ID>clock</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_DFF_LOW</type>
<position>72,-46</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>7 </output>
<input>
<ID>clock</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8</ID>
<type>AE_DFF_LOW</type>
<position>84,-46</position>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUT_0</ID>8 </output>
<input>
<ID>clock</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>42,-33</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>54,-33</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>66,-33</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>78,-33</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>52,-55</position>
<input>
<ID>N_in3</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>64,-55</position>
<input>
<ID>N_in3</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>76,-55</position>
<input>
<ID>N_in3</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>88,-55</position>
<input>
<ID>N_in3</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>CC_PULSE</type>
<position>39,-51</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-44,44.5,-33</points>
<intersection>-44 1</intersection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-44,45,-44</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>44,-33,44.5,-33</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-44,56.5,-33</points>
<intersection>-44 1</intersection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-44,57,-44</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-33,56.5,-33</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-44,68.5,-33</points>
<intersection>-44 1</intersection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-44,69,-44</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-33,68.5,-33</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-44,80.5,-33</points>
<intersection>-44 1</intersection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-44,81,-44</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80,-33,80.5,-33</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-54,52,-44</points>
<connection>
<GID>18</GID>
<name>N_in3</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-44,52,-44</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-54,64,-44</points>
<connection>
<GID>20</GID>
<name>N_in3</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-44,64,-44</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-54,76,-44</points>
<connection>
<GID>22</GID>
<name>N_in3</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-44,76,-44</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-54,88,-44</points>
<connection>
<GID>24</GID>
<name>N_in3</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-44,88,-44</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>88 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>45,-51,45,-47</points>
<connection>
<GID>2</GID>
<name>clock</name></connection>
<intersection>-51 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>41,-51,81,-51</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>45 3</intersection>
<intersection>57 6</intersection>
<intersection>69 8</intersection>
<intersection>81 10</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>57,-51,57,-47</points>
<connection>
<GID>4</GID>
<name>clock</name></connection>
<intersection>-51 4</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>69,-51,69,-47</points>
<connection>
<GID>6</GID>
<name>clock</name></connection>
<intersection>-51 4</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>81,-51,81,-47</points>
<connection>
<GID>8</GID>
<name>clock</name></connection>
<intersection>-51 4</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,182.7,-118</PageViewport></page 1>
<page 2>
<PageViewport>0,0,182.7,-118</PageViewport></page 2>
<page 3>
<PageViewport>0,0,182.7,-118</PageViewport></page 3>
<page 4>
<PageViewport>0,0,182.7,-118</PageViewport></page 4>
<page 5>
<PageViewport>0,0,182.7,-118</PageViewport></page 5>
<page 6>
<PageViewport>0,0,182.7,-118</PageViewport></page 6>
<page 7>
<PageViewport>0,0,182.7,-118</PageViewport></page 7>
<page 8>
<PageViewport>0,0,182.7,-118</PageViewport></page 8>
<page 9>
<PageViewport>0,0,182.7,-118</PageViewport></page 9></circuit>